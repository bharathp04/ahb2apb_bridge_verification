`ifndef ahb_apb_uvm_include_pkg
`define ahb_apb_uvm_include_pkg

package ahb_apb_uvm_include_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "ahb_apb_config.svh"
	`include "apb_slave_transaction.svh"
	`include "ahb_master_transaction.svh"
	`include "apb_slave_sequences.svh"
	`include "ahb_master_sequences.svh"
	`include "ahb_apb_virtual_sequences.svh"
	`include "apb_slave_sequencer.svh"
	`include "ahb_master_sequencer.svh"
	`include "ahb_master_driver.svh"
	`include "ahb_master_monitor.svh"
	`include "apb_slave_driver.svh"
	`include "apb_slave_monitor.svh"
	`include "ahb_master_agent.svh"
	`include "apb_slave_agent.svh"
	`include "ahb_apb_env.svh"
	`include "ahb_apb_tests.svh"
endpackage

import ahb_apb_uvm_include_pkg::*;

`endif