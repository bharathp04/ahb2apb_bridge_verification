package ahb_apb_bridge_pkg;
	parameter HADDR_SIZE= 32;
	parameter HDATA_SIZE= 32;
	
endpackage